library ieee;
use ieee.std_logic_1164.all;

package inst_pack is

constant nop1      : std_logic_vector( 5 downto 0) ;
constant xor1      : std_logic_vector( 5 downto 0) ;
constant and1      : std_logic_vector( 5 downto 0) ;
constant nxor1     : std_logic_vector( 5 downto 0) ;
constant nor1      : std_logic_vector( 5 downto 0) ;
constant nand1     : std_logic_vector( 5 downto 0) ;
constant add1      : std_logic_vector( 5 downto 0) ;
constant sub1      : std_logic_vector( 5 downto 0) ;
constant mul1      : std_logic_vector( 5 downto 0) ;
constant div1      : std_logic_vector( 5 downto 0) ;
constant addfp1    : std_logic_vector( 5 downto 0) ;
constant subfp1    : std_logic_vector( 5 downto 0) ;
constant mulfp1    : std_logic_vector( 5 downto 0) ;
constant divfp1    : std_logic_vector( 5 downto 0) ;
constant cmpreg1   : std_logic_vector( 5 downto 0) ;
constant not1      : std_logic_vector( 5 downto 0) ;
constant abs1      : std_logic_vector( 5 downto 0) ;
constant absfp1    : std_logic_vector( 5 downto 0) ;
constant sllr1     : std_logic_vector( 5 downto 0) ;
constant slar1     : std_logic_vector( 5 downto 0) ;
constant srlr1     : std_logic_vector( 5 downto 0) ;
constant srar1     : std_logic_vector( 5 downto 0) ;
constant rotlr1    : std_logic_vector( 5 downto 0) ;
constant rotrr1    : std_logic_vector( 5 downto 0) ;
constant ldr1      : std_logic_vector( 5 downto 0) ;
constant str1      : std_logic_vector( 5 downto 0) ;
constant xori1     : std_logic_vector( 5 downto 0) ;
constant andi1     : std_logic_vector( 5 downto 0) ;
constant ori1      : std_logic_vector( 5 downto 0) ;
constant nxori1    : std_logic_vector( 5 downto 0) ;
constant nori1     : std_logic_vector( 5 downto 0) ;
constant nandi1    : std_logic_vector( 5 downto 0) ;
constant addi1     : std_logic_vector( 5 downto 0) ;
constant subi1     : std_logic_vector( 5 downto 0) ;
constant muli1     : std_logic_vector( 5 downto 0) ;
constant divi1     : std_logic_vector( 5 downto 0) ;
constant addfpi1   : std_logic_vector( 5 downto 0) ;
constant subfpi1   : std_logic_vector( 5 downto 0) ;
constant mulfpi1   : std_logic_vector( 5 downto 0) ;
constant divfpi1   : std_logic_vector( 5 downto 0) ;
constant cmpregi1  : std_logic_vector( 5 downto 0) ;
constant jmp1      : std_logic_vector( 5 downto 0) ;
constant bre1      : std_logic_vector( 5 downto 0) ;
constant brue1     : std_logic_vector( 5 downto 0) ;
constant brg1      : std_logic_vector( 5 downto 0) ;
constant bls1      : std_logic_vector( 5 downto 0) ;
constant btr1      : std_logic_vector( 5 downto 0) ;
constant bfs1      : std_logic_vector( 5 downto 0) ;
constant jmpr1     : std_logic_vector( 5 downto 0) ; 
constant slli1     : std_logic_vector( 5 downto 0) ;
constant slai1     : std_logic_vector( 5 downto 0) ;
constant srli1     : std_logic_vector( 5 downto 0) ;
constant srai1     : std_logic_vector( 5 downto 0) ;
constant rotli1    : std_logic_vector( 5 downto 0) ;
constant rotri1    : std_logic_vector( 5 downto 0) ;
constant li1       : std_logic_vector( 5 downto 0) ;
constant ldm1      : std_logic_vector( 5 downto 0) ;
constant stm1      : std_logic_vector( 5 downto 0) ;
constant goto1     : std_logic_vector( 5 downto 0) ; 
constant mov1      : std_logic_vector( 5 downto 0) ;
constant clr1      : std_logic_vector( 5 downto 0) ;

constant R0   : std_logic_vector( 4 downto 0) ;
constant R1   : std_logic_vector( 4 downto 0) ;
constant R2   : std_logic_vector( 4 downto 0) ;
constant R3   : std_logic_vector( 4 downto 0) ;
constant R4   : std_logic_vector( 4 downto 0) ;
constant R5   : std_logic_vector( 4 downto 0) ;
constant R6   : std_logic_vector( 4 downto 0) ;
constant R7   : std_logic_vector( 4 downto 0) ;
constant R8   : std_logic_vector( 4 downto 0) ;
constant R9   : std_logic_vector( 4 downto 0) ;
constant R10  : std_logic_vector( 4 downto 0) ;
constant R11  : std_logic_vector( 4 downto 0) ;
constant R12  : std_logic_vector( 4 downto 0) ;
constant R13  : std_logic_vector( 4 downto 0) ;
constant R14  : std_logic_vector( 4 downto 0) ;
constant R15  : std_logic_vector( 4 downto 0) ;
constant R16  : std_logic_vector( 4 downto 0) ;
constant R17  : std_logic_vector( 4 downto 0) ;
constant R18  : std_logic_vector( 4 downto 0) ;
constant R19  : std_logic_vector( 4 downto 0) ;
constant R20  : std_logic_vector( 4 downto 0) ;
constant R21  : std_logic_vector( 4 downto 0) ;
constant R22  : std_logic_vector( 4 downto 0) ;
constant R23  : std_logic_vector( 4 downto 0) ;
constant R24  : std_logic_vector( 4 downto 0) ;
constant R25  : std_logic_vector( 4 downto 0) ;
constant R26  : std_logic_vector( 4 downto 0) ;
constant R27  : std_logic_vector( 4 downto 0) ;
constant R28  : std_logic_vector( 4 downto 0) ;
constant R29  : std_logic_vector( 4 downto 0) ;
constant R30  : std_logic_vector( 4 downto 0) ;
constant R31  : std_logic_vector( 4 downto 0) ;

end package inst_pack ;

package body inst_pack is

constant nop1      : std_logic_vector( 5 downto 0) :=  "000000" ;
constant xor1      : std_logic_vector( 5 downto 0) :=  "000001" ; 
constant and1      : std_logic_vector( 5 downto 0) :=  "000010" ;
constant nxor1     : std_logic_vector( 5 downto 0) :=  "000100" ;
constant nor1      : std_logic_vector( 5 downto 0) :=  "000101" ;
constant nand1     : std_logic_vector( 5 downto 0) :=  "000110" ;
constant add1      : std_logic_vector( 5 downto 0) :=  "000111" ;
constant sub1      : std_logic_vector( 5 downto 0) :=  "001000" ;
constant mul1      : std_logic_vector( 5 downto 0) :=  "001001" ;
constant div1      : std_logic_vector( 5 downto 0) :=  "001010" ;
constant addfp1    : std_logic_vector( 5 downto 0) :=  "001011" ;
constant subfp1    : std_logic_vector( 5 downto 0) :=  "001100" ;
constant mulfp1    : std_logic_vector( 5 downto 0) :=  "001101" ;
constant divfp1    : std_logic_vector( 5 downto 0) :=  "001110" ;
constant cmpreg1   : std_logic_vector( 5 downto 0) :=  "001111" ;
constant not1      : std_logic_vector( 5 downto 0) :=  "010000" ;
constant abs1      : std_logic_vector( 5 downto 0) :=  "010001" ;
constant absfp1    : std_logic_vector( 5 downto 0) :=  "010010" ;
constant sllr1     : std_logic_vector( 5 downto 0) :=  "010011" ;
constant slar1     : std_logic_vector( 5 downto 0) :=  "010100" ;
constant srlr1     : std_logic_vector( 5 downto 0) :=  "010101" ;
constant srar1     : std_logic_vector( 5 downto 0) :=  "010110" ;
constant rotlr1    : std_logic_vector( 5 downto 0) :=  "010111" ;
constant rotrr1    : std_logic_vector( 5 downto 0) :=  "011000" ;
constant ldr1      : std_logic_vector( 5 downto 0) :=  "011001" ;
constant str1      : std_logic_vector( 5 downto 0) :=  "011010" ;
constant xori1     : std_logic_vector( 5 downto 0) :=  "011011" ;
constant andi1     : std_logic_vector( 5 downto 0) :=  "011100" ;
constant ori1      : std_logic_vector( 5 downto 0) :=  "011101" ;
constant nxori1    : std_logic_vector( 5 downto 0) :=  "011110" ;
constant nori1     : std_logic_vector( 5 downto 0) :=  "011111" ;
constant nandi1    : std_logic_vector( 5 downto 0) :=  "100000" ;
constant addi1     : std_logic_vector( 5 downto 0) :=  "100001" ;
constant subi1     : std_logic_vector( 5 downto 0) :=  "100010" ;
constant muli1     : std_logic_vector( 5 downto 0) :=  "100011" ;
constant divi1     : std_logic_vector( 5 downto 0) :=  "100100" ;
constant addfpi1   : std_logic_vector( 5 downto 0) :=  "100101" ;
constant subfpi1   : std_logic_vector( 5 downto 0) :=  "100110" ;
constant mulfpi1   : std_logic_vector( 5 downto 0) :=  "100111" ;
constant divfpi1   : std_logic_vector( 5 downto 0) :=  "101000" ;
constant cmpregi1  : std_logic_vector( 5 downto 0) :=  "101001" ;
constant jmp1      : std_logic_vector( 5 downto 0) :=  "101010" ;
constant bre1      : std_logic_vector( 5 downto 0) :=  "101011" ;
constant brue1     : std_logic_vector( 5 downto 0) :=  "101100" ;
constant brg1      : std_logic_vector( 5 downto 0) :=  "101101" ;
constant bls1      : std_logic_vector( 5 downto 0) :=  "101110" ;
constant btr1      : std_logic_vector( 5 downto 0) :=  "101111" ;
constant bfs1      : std_logic_vector( 5 downto 0) :=  "110000" ;
constant jmpr1     : std_logic_vector( 5 downto 0) :=  "110001" ;
constant slli1     : std_logic_vector( 5 downto 0) :=  "110010" ;
constant slai1     : std_logic_vector( 5 downto 0) :=  "110011" ;
constant srli1     : std_logic_vector( 5 downto 0) :=  "110100" ;
constant srai1     : std_logic_vector( 5 downto 0) :=  "110101" ;
constant rotli1    : std_logic_vector( 5 downto 0) :=  "110110" ;
constant rotri1    : std_logic_vector( 5 downto 0) :=  "110111" ;
constant li1       : std_logic_vector( 5 downto 0) :=  "111000" ;
constant ldm1      : std_logic_vector( 5 downto 0) :=  "111001" ;
constant stm1      : std_logic_vector( 5 downto 0) :=  "111010" ;
constant goto1     : std_logic_vector( 5 downto 0) :=  "111111" ;
constant mov1      : std_logic_vector( 5 downto 0) :=  "111100" ;
constant clr1      : std_logic_vector( 5 downto 0) :=  "111101" ;

constant R0  : std_logic_vector( 4 downto 0)  :=  "00000" ;
constant R1  : std_logic_vector( 4 downto 0)  :=  "00001" ;
constant R2  : std_logic_vector( 4 downto 0)  :=  "00010" ;
constant R3  : std_logic_vector( 4 downto 0)  :=  "00011" ;
constant R4  : std_logic_vector( 4 downto 0)  :=  "00100" ;
constant R5  : std_logic_vector( 4 downto 0)  :=  "00101" ;
constant R6  : std_logic_vector( 4 downto 0)  :=  "00110" ;
constant R7  : std_logic_vector( 4 downto 0)  :=  "00111" ;
constant R8  : std_logic_vector( 4 downto 0)  :=  "01000" ;
constant R9  : std_logic_vector( 4 downto 0)  :=  "01001" ;
constant R10  : std_logic_vector( 4 downto 0) :=  "01010" ;
constant R11  : std_logic_vector( 4 downto 0) :=  "01011" ;
constant R12  : std_logic_vector( 4 downto 0) :=  "01100" ;
constant R13  : std_logic_vector( 4 downto 0) :=  "01101" ;
constant R14  : std_logic_vector( 4 downto 0) :=  "01110" ;
constant R15  : std_logic_vector( 4 downto 0) :=  "01111" ;
constant R16  : std_logic_vector( 4 downto 0) :=  "10000" ;
constant R17  : std_logic_vector( 4 downto 0) :=  "10001" ;
constant R18  : std_logic_vector( 4 downto 0) :=  "10010" ;
constant R19  : std_logic_vector( 4 downto 0) :=  "10011" ;
constant R20  : std_logic_vector( 4 downto 0) :=  "10100" ;
constant R21  : std_logic_vector( 4 downto 0) :=  "10101" ;
constant R22  : std_logic_vector( 4 downto 0) :=  "10110" ;
constant R23  : std_logic_vector( 4 downto 0) :=  "10111" ;
constant R24  : std_logic_vector( 4 downto 0) :=  "11000" ;
constant R25  : std_logic_vector( 4 downto 0) :=  "11001" ;
constant R26  : std_logic_vector( 4 downto 0) :=  "11010" ;
constant R27  : std_logic_vector( 4 downto 0) :=  "11011" ;
constant R28  : std_logic_vector( 4 downto 0) :=  "11100" ;
constant R29  : std_logic_vector( 4 downto 0) :=  "11101" ;
constant R30  : std_logic_vector( 4 downto 0) :=  "11110" ;
constant R31  : std_logic_vector( 4 downto 0) :=  "11111" ;

end package body inst_pack;



